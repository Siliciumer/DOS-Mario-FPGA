`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:         AGH UST
// Engineer: Wojciech Gredel, Hubert G�rowski
// 
// Create Date:    
// Design Name:     
// Module Name:     MarioFontRom
// Project Name:    DOS_Mario
// Target Devices:  Basys3
// Tool versions:   Vivado 2016.1
// Description:     
//	This module contains fonts
//  - 8-by-16 (8-by-2^4) font
//  - 20 characters (only necessary)
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - Module created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module MarioFontRom(
    input  wire [11:0] addr,            // {char_code[7:0], char_line[3:0]}
    output reg  [7:0]  char_line_pixels // pixels of the character line
    );

    // signal declaration
    reg [7:0] data;

    // body
    always @(*)
        char_line_pixels = data;

    always @*
        case (addr)
            //code x00
            12'h000: data = 8'b00000000; //
            12'h001: data = 8'b00000000; //  *****
            12'h002: data = 8'b01111100; // **   **
            12'h003: data = 8'b11000110; // **   **
            12'h004: data = 8'b11000110; // **  ***
            12'h005: data = 8'b11001110; // ** ****
            12'h006: data = 8'b11011110; // **** **
            12'h007: data = 8'b11110110; // ***  **
            12'h008: data = 8'b11100110; // **   **
            12'h009: data = 8'b11000110; // **   **
            12'h00a: data = 8'b11000110; //  *****
            12'h00b: data = 8'b01111100; //
            12'h00c: data = 8'b00000000; //
            12'h00d: data = 8'b00000000; //
            12'h00e: data = 8'b00000000; //
            12'h00f: data = 8'b00000000; //
            //code x01
            12'h010: data = 8'b00000000; //
            12'h011: data = 8'b00000000; //
            12'h012: data = 8'b00011000; //
            12'h013: data = 8'b00111000; //
            12'h014: data = 8'b01111000; //    **
            12'h015: data = 8'b00011000; //   ***
            12'h016: data = 8'b00011000; //  ****
            12'h017: data = 8'b00011000; //    **
            12'h018: data = 8'b00011000; //    **
            12'h019: data = 8'b00011000; //    **
            12'h01a: data = 8'b00011000; //    **
            12'h01b: data = 8'b00011000; //    **
            12'h01c: data = 8'b00011000; //    **
            12'h01d: data = 8'b00000000; //  ******
            12'h01e: data = 8'b00000000; //
            12'h01f: data = 8'b00000000; //
            //code x02
            12'h020: data = 8'b00000000; //
            12'h021: data = 8'b00000000; //
            12'h022: data = 8'b01111100; //  *****
            12'h023: data = 8'b11000110; // **   **
            12'h024: data = 8'b00000110; //      **
            12'h025: data = 8'b00001100; //     **
            12'h026: data = 8'b00011000; //    **
            12'h027: data = 8'b00110000; //   **
            12'h028: data = 8'b01100000; //  **
            12'h029: data = 8'b11000000; // **
            12'h02a: data = 8'b11000110; // **   **
            12'h02b: data = 8'b11111110; // *******
            12'h02c: data = 8'b00000000; //
            12'h02d: data = 8'b00000000; //
            12'h02e: data = 8'b00000000; //
            12'h02f: data = 8'b00000000; //
            //code x03
            12'h030: data = 8'b00000000; //
            12'h031: data = 8'b00000000; //
            12'h032: data = 8'b01111100; //  *****
            12'h033: data = 8'b11000110; // **   **
            12'h034: data = 8'b00000110; //      **
            12'h035: data = 8'b00000110; //      **
            12'h036: data = 8'b00111100; //   ****
            12'h037: data = 8'b00000110; //      **
            12'h038: data = 8'b00000110; //      **
            12'h039: data = 8'b00000110; //      **
            12'h03a: data = 8'b11000110; // **   **
            12'h03b: data = 8'b01111100; //  *****
            12'h03c: data = 8'b00000000; //
            12'h03d: data = 8'b00000000; //
            12'h03e: data = 8'b00000000; //
            12'h03f: data = 8'b00000000; //
            //code x04
            12'h040: data = 8'b00000000; //
            12'h041: data = 8'b00000000; //
            12'h042: data = 8'b00001100; //     **
            12'h043: data = 8'b00011100; //    ***
            12'h044: data = 8'b00111100; //   ****
            12'h045: data = 8'b01101100; //  ** **
            12'h046: data = 8'b11001100; // **  **
            12'h047: data = 8'b11111110; // *******
            12'h048: data = 8'b00001100; //     **
            12'h049: data = 8'b00001100; //     **
            12'h04a: data = 8'b00001100; //     **
            12'h04b: data = 8'b00011110; //    ****
            12'h04c: data = 8'b00000000; //
            12'h04d: data = 8'b00000000; //
            12'h04e: data = 8'b00000000; //
            12'h04f: data = 8'b00000000; //
            //code x05
            12'h050: data = 8'b00000000; //
            12'h051: data = 8'b00000000; //
            12'h052: data = 8'b11111110; // *******
            12'h053: data = 8'b11000000; // **
            12'h054: data = 8'b11000000; // **
            12'h055: data = 8'b11000000; // **
            12'h056: data = 8'b11111100; // ******
            12'h057: data = 8'b00000110; //      **
            12'h058: data = 8'b00000110; //      **
            12'h059: data = 8'b00000110; //      **
            12'h05a: data = 8'b11000110; // **   **
            12'h05b: data = 8'b01111100; //  *****
            12'h05c: data = 8'b00000000; //
            12'h05d: data = 8'b00000000; //
            12'h05e: data = 8'b00000000; //
            12'h05f: data = 8'b00000000; //
            //code x06
            12'h060: data = 8'b00000000; //
            12'h061: data = 8'b00000000; //
            12'h062: data = 8'b00111000; //   ***
            12'h063: data = 8'b01100000; //  **
            12'h064: data = 8'b11000000; // **
            12'h065: data = 8'b11000000; // **
            12'h066: data = 8'b11111100; // ******
            12'h067: data = 8'b11000110; // **   **
            12'h068: data = 8'b11000110; // **   **
            12'h069: data = 8'b11000110; // **   **
            12'h06a: data = 8'b11000110; // **   **
            12'h06b: data = 8'b01111100; //  *****
            12'h06c: data = 8'b00000000; //
            12'h06d: data = 8'b00000000; //
            12'h06e: data = 8'b00000000; //
            12'h06f: data = 8'b00000000; //
            //code x07
            12'h070: data = 8'b00000000; //
            12'h071: data = 8'b00000000; //
            12'h072: data = 8'b11111110; // *******
            12'h073: data = 8'b11000110; // **   **
            12'h074: data = 8'b00000110; //      **
            12'h075: data = 8'b00000110; //      **
            12'h076: data = 8'b00001100; //     **
            12'h077: data = 8'b00011000; //    **
            12'h078: data = 8'b00110000; //   **
            12'h079: data = 8'b00110000; //   **
            12'h07a: data = 8'b00110000; //   **
            12'h07b: data = 8'b00110000; //   **
            12'h07c: data = 8'b00000000; //
            12'h07d: data = 8'b00000000; //
            12'h07e: data = 8'b00000000; //
            12'h07f: data = 8'b00000000; //
            //code x08
            12'h080: data = 8'b00000000; //
            12'h081: data = 8'b00000000; //
            12'h082: data = 8'b01111100; //  *****
            12'h083: data = 8'b11000110; // **   **
            12'h084: data = 8'b11000110; // **   **
            12'h085: data = 8'b11000110; // **   **
            12'h086: data = 8'b01111100; //  *****
            12'h087: data = 8'b11000110; // **   **
            12'h088: data = 8'b11000110; // **   **
            12'h089: data = 8'b11000110; // **   **
            12'h08a: data = 8'b11000110; // **   **
            12'h08b: data = 8'b01111100; //  *****
            12'h08c: data = 8'b00000000; //
            12'h08d: data = 8'b00000000; //
            12'h08e: data = 8'b00000000; //
            12'h08f: data = 8'b00000000; //
            //code x09
            12'h090: data = 8'b00000000; //
            12'h091: data = 8'b00000000; //
            12'h092: data = 8'b01111100; //  *****
            12'h093: data = 8'b11000110; // **   **
            12'h094: data = 8'b11000110; // **   **
            12'h095: data = 8'b11000110; // **   **
            12'h096: data = 8'b01111110; //  ******
            12'h097: data = 8'b00000110; //      **
            12'h098: data = 8'b00000110; //      **
            12'h099: data = 8'b00000110; //      **
            12'h09a: data = 8'b00001100; //     **
            12'h09b: data = 8'b01111000; //  ****
            12'h09c: data = 8'b00000000; //
            12'h09d: data = 8'b00000000; //
            12'h09e: data = 8'b00000000; //
            12'h09f: data = 8'b00000000; //
            //code x0a
            12'h0a0: data = 8'b00000000; //
            12'h0a1: data = 8'b00000000; //
            12'h0a2: data = 8'b11000011; // **    **
            12'h0a3: data = 8'b11100111; // ***  ***
            12'h0a4: data = 8'b11111111; // ********
            12'h0a5: data = 8'b11111111; // ********
            12'h0a6: data = 8'b11011011; // ** ** **
            12'h0a7: data = 8'b11000011; // **    **
            12'h0a8: data = 8'b11000011; // **    **
            12'h0a9: data = 8'b11000011; // **    **
            12'h0aa: data = 8'b11000011; // **    **
            12'h0ab: data = 8'b11000011; // **    **
            12'h0ac: data = 8'b00000000; //
            12'h0ad: data = 8'b00000000; //
            12'h0ae: data = 8'b00000000; //
            12'h0af: data = 8'b00000000; //
            //code x0b
            12'h0b0: data = 8'b00000000; //
            12'h0b1: data = 8'b00000000; //
            12'h0b2: data = 8'b00010000; //    *
            12'h0b3: data = 8'b00111000; //   ***
            12'h0b4: data = 8'b01101100; //  ** **
            12'h0b5: data = 8'b11000110; // **   **
            12'h0b6: data = 8'b11000110; // **   **
            12'h0b7: data = 8'b11111110; // *******
            12'h0b8: data = 8'b11000110; // **   **
            12'h0b9: data = 8'b11000110; // **   **
            12'h0ba: data = 8'b11000110; // **   **
            12'h0bb: data = 8'b11000110; // **   **
            12'h0bc: data = 8'b00000000; //
            12'h0bd: data = 8'b00000000; //
            12'h0be: data = 8'b00000000; //
            12'h0bf: data = 8'b00000000; //
            //code x0c
            12'h0c0: data = 8'b00000000; //
            12'h0c1: data = 8'b00000000; //
            12'h0c2: data = 8'b11111100; // ******
            12'h0c3: data = 8'b01100110; //  **  **
            12'h0c4: data = 8'b01100110; //  **  **
            12'h0c5: data = 8'b01100110; //  **  **
            12'h0c6: data = 8'b01111100; //  *****
            12'h0c7: data = 8'b01101100; //  ** **
            12'h0c8: data = 8'b01100110; //  **  **
            12'h0c9: data = 8'b01100110; //  **  **
            12'h0ca: data = 8'b01100110; //  **  **
            12'h0cb: data = 8'b11100110; // ***  **
            12'h0cc: data = 8'b00000000; //
            12'h0cd: data = 8'b00000000; //
            12'h0ce: data = 8'b00000000; //
            12'h0cf: data = 8'b00000000; //
            //code x0d
            12'h0d0: data = 8'b00000000; //
            12'h0d1: data = 8'b00000000; //
            12'h0d2: data = 8'b00111100; //   ****
            12'h0d3: data = 8'b00011000; //    **
            12'h0d4: data = 8'b00011000; //    **
            12'h0d5: data = 8'b00011000; //    **
            12'h0d6: data = 8'b00011000; //    **
            12'h0d7: data = 8'b00011000; //    **
            12'h0d8: data = 8'b00011000; //    **
            12'h0d9: data = 8'b00011000; //    **
            12'h0da: data = 8'b00011000; //    **
            12'h0db: data = 8'b00111100; //   ****
            12'h0dc: data = 8'b00000000; //
            12'h0dd: data = 8'b00000000; //
            12'h0de: data = 8'b00000000; //
            12'h0df: data = 8'b00000000; //
            //code x0e
            12'h0e0: data = 8'b00000000; //
            12'h0e1: data = 8'b00000000; //
            12'h0e2: data = 8'b01111100; //  *****
            12'h0e3: data = 8'b11000110; // **   **
            12'h0e4: data = 8'b11000110; // **   **
            12'h0e5: data = 8'b11000110; // **   **
            12'h0e6: data = 8'b11000110; // **   **
            12'h0e7: data = 8'b11000110; // **   **
            12'h0e8: data = 8'b11000110; // **   **
            12'h0e9: data = 8'b11000110; // **   **
            12'h0ea: data = 8'b11000110; // **   **
            12'h0eb: data = 8'b01111100; //  *****
            12'h0ec: data = 8'b00000000; //
            12'h0ed: data = 8'b00000000; //
            12'h0ee: data = 8'b00000000; //
            12'h0ef: data = 8'b00000000; //
            //code x0f
            12'h0f0: data = 8'b00000000; //
            12'h0f1: data = 8'b00000000; //
            12'h0f2: data = 8'b00000000; //
            12'h0f3: data = 8'b00000000; //
            12'h0f4: data = 8'b00000000; //
            12'h0f5: data = 8'b00000000; //
            12'h0f6: data = 8'b00000000; //
            12'h0f7: data = 8'b00000000; //
            12'h0f8: data = 8'b00000000; //
            12'h0f9: data = 8'b00000000; //
            12'h0fa: data = 8'b00000000; //
            12'h0fb: data = 8'b00000000; //
            12'h0fc: data = 8'b00000000; //
            12'h0fd: data = 8'b00000000; //
            12'h0fe: data = 8'b00000000; //
            12'h0ff: data = 8'b00000000; //
            //code x10
            12'h100: data = 8'b00000000; //
            12'h101: data = 8'b00000000; //
            12'h102: data = 8'b00000000; //
            12'h103: data = 8'b00000000; //
            12'h104: data = 8'b00000000; //
            12'h105: data = 8'b11000011; // **    **
            12'h106: data = 8'b01100110; //  **  **
            12'h107: data = 8'b00111100; //   ****
            12'h108: data = 8'b00011000; //    **
            12'h109: data = 8'b00111100; //   ****
            12'h10a: data = 8'b01100110; //  **  **
            12'h10b: data = 8'b11000011; // **    **
            12'h10c: data = 8'b00000000; //
            12'h10d: data = 8'b00000000; //
            12'h10e: data = 8'b00000000; //
            12'h10f: data = 8'b00000000; //
            //code x11
            12'h110: data = 8'b00000000; //
            12'h111: data = 8'b00000000; //
            12'h112: data = 8'b00000000; //
            12'h113: data = 8'b00000000; //  
            12'h114: data = 8'b00111100; //   ****
            12'h115: data = 8'b00111100; //   ****
            12'h116: data = 8'b11111111; // **    **
            12'h117: data = 8'b11111111; // **    **
            12'h118: data = 8'b11111111; // **    **
            12'h119: data = 8'b11111111; // **    **
            12'h11a: data = 8'b00111100; //   ****
            12'h11b: data = 8'b00111100; //   ****
            12'h11c: data = 8'b00000000; //
            12'h11d: data = 8'b00000000; //
            12'h11e: data = 8'b00000000; //
            12'h11f: data = 8'b00000000; //
            //code x12
            12'h120: data = 8'b00000000; //
            12'h121: data = 8'b00000000; //
            12'h122: data = 8'b11110000; // ****
            12'h123: data = 8'b01100000; //  **
            12'h124: data = 8'b01100000; //  **
            12'h125: data = 8'b01100000; //  **
            12'h126: data = 8'b01100000; //  **
            12'h127: data = 8'b01100000; //  **
            12'h128: data = 8'b01100000; //  **
            12'h129: data = 8'b01100010; //  **   *
            12'h12a: data = 8'b01100110; //  **  **
            12'h12b: data = 8'b11111110; // *******
            12'h12c: data = 8'b00000000; //
            12'h12d: data = 8'b00000000; //
            12'h12e: data = 8'b00000000; //
            12'h12f: data = 8'b00000000; //
            //code x13
            12'h130: data = 8'b00000000; //
            12'h131: data = 8'b00000000; //
            12'h132: data = 8'b11111110; // *******
            12'h133: data = 8'b01100110; //  **  **
            12'h134: data = 8'b01100010; //  **   *
            12'h135: data = 8'b01101000; //  ** *
            12'h136: data = 8'b01111000; //  ****
            12'h137: data = 8'b01111000; //  ****
            12'h138: data = 8'b01101000; //  ** *
            12'h139: data = 8'b01100010; //  **   *
            12'h13a: data = 8'b01100110; //  **  **
            12'h13b: data = 8'b11111110; // *******
            12'h13c: data = 8'b00000000; //
            12'h13d: data = 8'b00000000; //
            12'h13e: data = 8'b00000000; //
            12'h13f: data = 8'b00000000; //
            //code x14
            12'h140: data = 8'b00000000; //
            12'h141: data = 8'b00000000; //
            12'h142: data = 8'b11000011; // **    **
            12'h143: data = 8'b11000011; // **    **
            12'h144: data = 8'b11000011; // **    **
            12'h145: data = 8'b11000011; // **    **
            12'h146: data = 8'b11000011; // **    **
            12'h147: data = 8'b11000011; // **    **
            12'h148: data = 8'b11000011; // **    **
            12'h149: data = 8'b01100110; //  **  **
            12'h14a: data = 8'b00111100; //   ****
            12'h14b: data = 8'b00011000; //    **
            12'h14c: data = 8'b00000000; //
            12'h14d: data = 8'b00000000; //
            12'h14e: data = 8'b00000000; //
            12'h14f: data = 8'b00000000; //
            
            default: data = 8'b00000000;
        endcase

endmodule
